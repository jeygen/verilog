// Avoid metastability from fast to slow clocks
// 
