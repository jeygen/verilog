new module pattern_detect(
