wire a [5-1:0]
// is equiv to
wire a [4:0]

// if integer than vector is elements not bits, prob be 32 bits each
integer a [4:0]

// order is a style issue
wire [3:0] b;
wire b [3:0];
