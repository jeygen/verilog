// program dual ff synchronizer fast to slow, and slow to fast
// program RAM
