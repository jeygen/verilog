// code a alu with modules
