two types of asserts: immediate and concurrent

concurrent use "assert property"
if condition is true nothing happens
  'disable iff' allows conditional skipping of assert property
