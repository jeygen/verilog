bit: A binary digit that can have one of two values: 0 or 1.
byte: An 8-bit data type.
shortint: A signed 16-bit integer.
int: A signed 32-bit integer.
longint: A signed 64-bit integer.
real: A single-precision floating-point number.
realtime: A double-precision floating-point number.
logic: A four-state data type that can have one of four values: 0, 1, X (unknown), or Z (high impedance).
reg: A one-bit or multi-bit data type that can be used to represent a register, think more "evaluated at a certian point"
automatic: This qualifier means created and destroyed with function among other things, for non-static things
