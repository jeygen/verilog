// do this
