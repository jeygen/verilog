// Practice Here

