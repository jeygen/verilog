// fpga embedded ram = block ram
// max bram diff for diff fpga
// width x depth = size
// diff configs avail: single, dual. fifo
