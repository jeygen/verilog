// Practice Here
