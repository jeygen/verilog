// Avoid metastability when going from slow to fast
