// lets go

	

