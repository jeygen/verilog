// for crossing domains when more than just a pulse
