/*

Levels of verilog abstraction: 
  Behavioral level:
    Concurrent algos. Each algo is sequential, consists of set of instrucitons
    executed in sequence. Functions, Tasks, Always blocks. No regard for structure.
  Register-Transfer Level:
    RTL is data b/t reg. Explicit clk used. Exact timing. Anything sythesizable is RTL.
  Gate Level:	
    Within the logic level the characteristics of a system are described by logical links and their timing properties. 
    All signals are discrete signals. They can only have definite logical values (`0', `1', `X', `Z`). 
    The usable operations are predefined logic primitives (AND, OR, NOT etc gates). Using gate level modeling might not be a good idea for any level of logic design. 
    Gate level code is generated by tools like synthesis tools and this netlist is used for gate level simulation and for backend.
    
  This tut:
    Specifications (specs)
    High level design
    Low level (micro) design
    RTL coding
    Verification
    Synthesis.
    
 */
