/*
initial can be used instead of always
both execute a sim from timecode 0 and go to end of block but inital just happens once
*/
